
module instr_mem(
    input [31:0] addr,
    output logic [31:0] instr
    );
    logic [31:0] mem [1023:0];
/*    
    initial begin
        mem[0] = 32'b00000000001000001000000110110011; //ADD x3, x1, x2
        mem[1] = 32'b0100000_00100_00011_000_00110_0110011; //SUB x6, x3, x4
        mem[2] = 32'b00000000111100111111010000010011; //ANDI x8, x7, 15
        mem[3] = 32'b00000000101000010010010010010011; //SLTI x9, x2, 10
        mem[4] = 32'b00000000010100111010010100000011; //LW x10, 5(x7)
        mem[5] = 32'b11111111110000010010010110000011; //LW x11, -4(x2)
        mem[6] = 32'b00000000000100100010010100100011; //SW x1, 10(x4)
        mem[7] = 32'b11111110010100010010111110100011; //SW x5, -1(x2)
        mem[8] = 32'b00000000110000001101010001100011; //BGE x1, x12, 8
        mem[9] = 32'b00000000001000001001011010110011; //SLL x13, x1, x2
        mem[10] = 32'b00000000001000001101011010110011; //SRL x13, x1, x2
        mem[11] = 32'b00010010001101000101011100110111; //LUI x14, 0x12345            
        mem[12] = 32'b01100111100010010000011110010111; //AUIPC x15, 0x67890
        mem[13] = 32'b0_0001000000_0_00000000_11010_1101111; //JAL x26, 128
        mem[45] = 32'b00000000000011010000110111100111; //JALR x27, x26, 0
    end
 */   
    
    /*
    initial begin
        $readmemh("C:\\Users\\HP\\Desktop\\tb_6\\instr.txt",mem);
    end
    */
    
    assign instr = mem[addr >> 2];
endmodule

