
module Add(
    input logic [31:0] operand1,operand2,
    output logic [31:0] result
    );
    assign  result = operand1 + operand2;
endmodule

