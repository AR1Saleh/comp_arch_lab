
module PC_Adder(
    input logic [31:0] operand1,
    output logic [31:0] result
    );
    assign  result = operand1 + 4;
endmodule

